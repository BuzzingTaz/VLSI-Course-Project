* SPICE3 file created from or.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY=1.8
.option scale=0.09u
.global vdd gnd

Vdd vdd gnd SUPPLY
Va A gnd pulse 0 1.8 0ns 0.1ns 0.1ns 9.9ns 20ns
Vb B gnd pulse 0 1.8 0ns 0.1ns 0.1ns 19.9ns 40ns

M1000 orout a_13_n15# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=60 ps=54
M1001 a_13_n15# B a_13_9# w_0_3# CMOSP w=8 l=2
+  ad=40 pd=26 as=64 ps=32
M1002 gnd B a_13_n15# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1003 a_13_9# A vdd w_0_3# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=52
M1004 a_13_n15# A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 orout a_13_n15# vdd w_0_3# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
.tran 0.1n 80n

.control
run
plot v(A)
plot v(B)

plot  v(orout)

.endc
.end