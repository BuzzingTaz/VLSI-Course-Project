magic
tech scmos
timestamp 1638828401
<< metal1 >>
rect -10 324 102 328
rect 180 324 546 328
rect 11 300 101 304
rect 176 300 181 304
rect 196 300 227 304
rect 286 300 290 304
rect 304 300 329 304
rect 396 300 405 304
rect 450 300 482 304
rect 20 293 101 297
rect 205 293 227 297
rect 313 293 331 297
rect 405 293 406 297
rect 456 293 482 297
rect 563 293 565 297
rect 29 286 101 290
rect 214 286 227 290
rect 322 286 334 290
rect 465 286 483 290
rect 38 279 101 283
rect 223 279 231 283
rect 474 279 483 283
rect 47 272 100 276
rect 404 275 408 278
rect 384 271 408 275
rect 322 268 326 271
rect 189 264 227 268
rect 293 264 326 268
rect 450 268 454 278
rect 450 264 485 268
rect 189 261 192 264
rect 482 261 485 264
rect -1 257 103 261
rect 181 257 192 261
rect 386 256 450 260
rect 295 249 459 253
rect 186 241 468 245
rect 29 233 190 237
rect 38 225 199 229
rect 204 225 298 229
rect 47 217 208 221
rect 213 217 307 221
rect 312 217 390 221
rect 55 209 218 213
rect 64 202 316 206
rect 73 195 399 199
rect 82 188 479 192
rect -31 180 -15 184
rect -10 180 421 184
rect 11 156 106 160
rect 165 156 169 160
rect 183 156 208 160
rect 275 156 284 160
rect 329 156 357 160
rect 421 156 424 160
rect 20 149 106 153
rect 192 149 210 153
rect 284 149 285 153
rect 335 149 356 153
rect 29 142 106 146
rect 201 142 213 146
rect 344 142 356 146
rect 38 135 110 139
rect 283 131 287 134
rect 263 127 287 131
rect 201 124 205 127
rect -27 120 -6 124
rect -1 120 106 124
rect 172 120 205 124
rect 329 124 333 134
rect 329 120 357 124
rect 265 112 329 116
rect 174 105 338 109
rect 29 96 177 100
rect 38 88 186 92
rect 191 88 269 92
rect 55 80 195 84
rect 64 72 278 76
rect 73 64 347 68
rect -10 55 251 59
rect 11 31 101 35
rect 155 31 159 35
rect 173 31 183 35
rect 227 31 248 35
rect 20 24 100 28
rect 182 24 184 28
rect 222 27 223 31
rect 239 24 248 28
rect 308 21 311 25
rect 29 17 103 21
rect 179 6 182 9
rect -1 2 182 6
rect 226 6 229 9
rect 226 2 252 6
rect -41 -13 5 -9
rect 10 -13 329 -9
rect -41 -27 15 -23
rect 164 -24 233 -20
rect -41 -35 24 -31
rect 29 -35 167 -31
rect -41 -43 32 -39
rect -41 -51 41 -47
rect -41 -60 50 -56
rect 55 -60 176 -56
rect -41 -69 58 -65
rect 63 -69 242 -65
rect -41 -78 67 -74
rect -41 -85 76 -81
rect 55 -93 155 -89
rect -10 -101 191 -97
rect 20 -125 107 -121
rect 150 -125 174 -121
rect 215 -125 218 -121
rect 10 -132 117 -128
rect 160 -132 173 -128
rect -2 -147 191 -143
<< m2contact >>
rect -15 323 -10 328
rect 6 299 11 304
rect 181 299 186 304
rect 191 299 196 304
rect 290 299 295 304
rect 299 299 304 304
rect 381 299 386 304
rect 391 299 396 304
rect 15 292 20 297
rect 200 292 205 297
rect 308 292 313 297
rect 400 292 405 297
rect 451 292 456 297
rect 24 285 29 290
rect 209 285 214 290
rect 317 285 322 290
rect 460 285 465 290
rect 33 278 38 283
rect 218 278 223 283
rect 469 278 474 283
rect 42 271 47 276
rect 478 271 483 276
rect -6 256 -1 261
rect 381 256 386 261
rect 450 256 455 261
rect 290 249 295 254
rect 459 249 464 254
rect 181 241 186 246
rect 468 241 473 246
rect 24 233 29 238
rect 190 233 195 238
rect 33 225 38 230
rect 199 225 204 230
rect 298 225 303 230
rect 42 217 47 222
rect 208 217 213 222
rect 307 217 312 222
rect 390 217 395 222
rect 50 208 55 213
rect 218 209 223 214
rect 59 201 64 206
rect 316 202 321 207
rect 68 194 73 199
rect 399 195 404 200
rect 77 187 82 192
rect 479 188 484 193
rect -15 179 -10 184
rect 6 155 11 160
rect 169 155 174 160
rect 178 155 183 160
rect 260 155 265 160
rect 270 155 275 160
rect 15 148 20 153
rect 187 148 192 153
rect 279 148 284 153
rect 330 148 335 153
rect 24 141 29 146
rect 196 141 201 146
rect 339 141 344 146
rect 33 134 38 139
rect 348 134 353 139
rect -6 119 -1 124
rect 260 112 265 117
rect 329 112 334 117
rect 169 105 174 110
rect 338 104 343 109
rect 24 96 29 101
rect 177 96 182 101
rect 33 88 38 93
rect 186 88 191 93
rect 269 88 274 93
rect 50 80 55 85
rect 195 80 200 85
rect 59 71 64 76
rect 278 72 283 77
rect 68 63 73 68
rect 347 64 352 69
rect -15 55 -10 60
rect 6 30 11 35
rect 159 30 164 35
rect 168 30 173 35
rect 15 23 20 28
rect 177 23 182 28
rect 234 23 239 28
rect 24 16 29 21
rect 243 16 248 21
rect -6 2 -1 7
rect 5 -14 10 -9
rect 15 -27 20 -22
rect 159 -25 164 -20
rect 233 -24 238 -19
rect 24 -35 29 -30
rect 167 -35 172 -30
rect 32 -44 37 -39
rect 41 -51 46 -46
rect 50 -60 55 -55
rect 176 -60 181 -55
rect 58 -70 63 -65
rect 242 -69 247 -64
rect 67 -78 72 -73
rect 76 -85 81 -80
rect 50 -93 55 -88
rect 155 -94 160 -89
rect -15 -101 -10 -96
rect 15 -125 20 -120
rect 5 -133 10 -128
rect 155 -133 160 -128
rect -7 -147 -2 -142
<< metal2 >>
rect -15 184 -11 323
rect -15 60 -11 179
rect -6 124 -2 256
rect 6 160 10 299
rect -15 -96 -11 55
rect -6 7 -2 119
rect 6 35 10 155
rect 15 153 19 292
rect 24 238 28 285
rect -6 -142 -2 2
rect 6 -9 10 30
rect 6 -128 10 -14
rect 15 28 19 148
rect 24 146 28 233
rect 33 230 37 278
rect 24 101 28 141
rect 33 139 37 225
rect 42 222 46 271
rect 181 246 185 299
rect 191 238 195 299
rect 200 230 204 292
rect 209 222 213 285
rect 15 -22 19 23
rect 24 21 28 96
rect 33 93 37 134
rect 15 -120 19 -27
rect 24 -30 28 16
rect 33 -39 37 88
rect 42 -46 46 217
rect 218 214 222 278
rect 291 254 295 299
rect 299 230 303 299
rect 308 222 312 292
rect 50 85 54 208
rect 317 207 321 285
rect 382 261 386 299
rect 391 222 395 299
rect 50 -55 54 80
rect 59 76 63 201
rect 400 200 404 292
rect 451 261 455 292
rect 460 254 464 285
rect 469 246 473 278
rect 50 -88 54 -60
rect 59 -65 63 71
rect 68 68 72 194
rect 478 193 482 271
rect 68 -73 72 63
rect 77 -80 81 187
rect 170 110 174 155
rect 178 101 182 155
rect 187 93 191 148
rect 196 85 200 141
rect 261 117 265 155
rect 270 93 274 155
rect 279 77 283 148
rect 330 117 334 148
rect 339 109 343 141
rect 348 69 352 134
rect 160 -20 164 30
rect 168 -30 172 30
rect 177 -55 181 23
rect 234 -19 238 23
rect 243 -64 247 16
rect 156 -128 160 -94
use and5  and5_0
timestamp 1638797340
transform 1 0 100 0 1 304
box 0 -47 82 24
use and4  and4_1
timestamp 1638631971
transform 1 0 221 0 1 304
box 0 -40 72 24
use and3  and3_2
timestamp 1638770576
transform 1 0 322 0 1 304
box 0 -33 62 24
use and  and_3
timestamp 1638780161
transform 1 0 404 0 1 301
box 0 -23 50 27
use or5  or5_0
timestamp 1638800402
transform 1 0 482 0 1 301
box 0 -44 81 27
use and4  and4_0
timestamp 1638631971
transform 1 0 100 0 1 160
box 0 -40 72 24
use and3  and3_1
timestamp 1638770576
transform 1 0 201 0 1 160
box 0 -33 62 24
use and  and_2
timestamp 1638780161
transform 1 0 283 0 1 157
box 0 -23 50 27
use or4  or4_0
timestamp 1638782314
transform 1 0 350 0 1 157
box 0 -37 71 27
use and3  and3_0
timestamp 1638770576
transform 1 0 100 0 1 35
box 0 -33 62 24
use and  and_1
timestamp 1638780161
transform 1 0 179 0 1 32
box 0 -23 50 27
use or3  or3_0
timestamp 1638771050
transform 1 0 247 0 1 32
box 0 -30 61 27
use and  and_0
timestamp 1638780161
transform 1 0 100 0 1 -124
box 0 -23 50 27
use or  or_0
timestamp 1638780148
transform 1 0 165 0 1 -124
box 0 -23 50 27
<< labels >>
rlabel metal1 -31 180 -29 184 5 vdd
rlabel metal1 -27 120 -25 124 1 gnd
rlabel metal1 421 156 424 160 7 C3
rlabel metal1 308 21 311 25 1 C2
rlabel metal1 564 295 564 295 7 C4
rlabel metal1 -41 -78 -38 -74 3 G2
rlabel metal1 -41 -85 -38 -81 3 G3
rlabel metal1 -41 -69 -38 -65 3 G1
rlabel metal1 -41 -60 -38 -56 3 G0
rlabel metal1 -41 -51 -38 -47 3 P3
rlabel metal1 -41 -43 -38 -39 3 P2
rlabel metal1 -41 -35 -38 -31 3 P1
rlabel metal1 -41 -27 -38 -23 3 P0
rlabel metal1 215 -125 218 -121 1 C1
rlabel metal1 -41 -13 -38 -9 3 C0
<< end >>
