magic
tech scmos
timestamp 1638631971
<< nwell >>
rect 0 0 72 20
<< ntransistor >>
rect 12 -32 14 -28
rect 22 -32 24 -28
rect 32 -32 34 -28
rect 42 -32 44 -28
rect 59 -32 61 -28
<< ptransistor >>
rect 12 6 14 14
rect 22 6 24 14
rect 32 6 34 14
rect 42 6 44 14
rect 59 6 61 14
<< ndiffusion >>
rect 10 -32 12 -28
rect 14 -32 22 -28
rect 24 -32 32 -28
rect 34 -32 42 -28
rect 44 -32 46 -28
rect 58 -32 59 -28
rect 61 -32 62 -28
<< pdiffusion >>
rect 10 6 12 14
rect 14 6 16 14
rect 20 6 22 14
rect 24 6 26 14
rect 30 6 32 14
rect 34 6 36 14
rect 40 6 42 14
rect 44 6 46 14
rect 58 6 59 14
rect 61 6 62 14
<< ndcontact >>
rect 6 -32 10 -28
rect 46 -32 50 -28
rect 54 -32 58 -28
rect 62 -32 66 -28
<< pdcontact >>
rect 6 6 10 14
rect 16 6 20 14
rect 26 6 30 14
rect 36 6 40 14
rect 46 6 50 14
rect 54 6 58 14
rect 62 6 66 14
<< polysilicon >>
rect 12 14 14 17
rect 22 14 24 17
rect 32 14 34 17
rect 42 14 44 17
rect 59 14 61 17
rect 12 -28 14 6
rect 22 -28 24 6
rect 32 -28 34 6
rect 42 -28 44 6
rect 59 -28 61 6
rect 12 -35 14 -32
rect 22 -35 24 -32
rect 32 -35 34 -32
rect 42 -35 44 -32
rect 59 -35 61 -32
<< polycontact >>
rect 8 -4 12 0
rect 18 -11 22 -7
rect 28 -18 32 -14
rect 38 -25 42 -21
rect 55 -4 59 0
<< metal1 >>
rect 0 20 72 24
rect 6 14 10 20
rect 26 14 30 20
rect 46 14 50 20
rect 54 14 58 20
rect 16 0 20 6
rect 36 0 40 6
rect 62 0 66 6
rect 0 -4 8 0
rect 16 -4 55 0
rect 62 -4 72 0
rect 0 -11 18 -7
rect 0 -18 28 -14
rect 0 -25 38 -21
rect 46 -28 50 -4
rect 62 -28 66 -4
rect 6 -36 10 -32
rect 54 -36 58 -32
rect 0 -40 72 -36
<< labels >>
rlabel metal1 1 -2 1 -2 3 A
rlabel metal1 1 -9 1 -9 3 B
rlabel metal1 2 22 2 22 4 vdd
rlabel metal1 2 -38 2 -38 2 gnd
rlabel metal1 1 -23 1 -23 3 D
rlabel metal1 70 -2 70 -2 7 out
rlabel metal1 1 -16 1 -16 3 C
<< end >>
