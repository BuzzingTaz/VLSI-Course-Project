magic
tech scmos
timestamp 1638828310
<< metal1 >>
rect 1172 382 1230 386
rect 1177 351 1220 355
rect 495 238 583 242
rect 495 169 499 238
rect 1037 214 1213 218
rect 510 178 586 182
rect 485 165 499 169
rect 924 82 1206 83
rect 921 79 1206 82
rect 917 59 921 64
rect 498 45 576 49
rect 572 43 576 45
rect 498 31 544 35
rect 549 31 576 35
rect 1202 31 1206 79
rect 1209 39 1213 214
rect 1216 47 1220 351
rect 1226 137 1230 382
rect 1739 119 1743 123
rect 1739 111 1743 115
rect 1739 103 1743 107
rect 1739 91 1743 95
rect 1216 43 1230 47
rect 1209 35 1232 39
rect 497 23 535 27
rect 1202 27 1227 31
rect 540 23 575 27
rect 499 15 526 19
rect 1187 19 1230 23
rect 531 15 577 19
rect 499 7 517 11
rect 522 7 577 11
rect 486 -2 576 2
rect 483 -11 576 -7
rect 484 -20 577 -16
rect 485 -27 578 -23
rect 496 -49 504 -45
rect 1187 -63 1191 19
rect 828 -66 1191 -63
rect 831 -67 1191 -66
rect 1194 6 1234 10
rect 1194 -93 1198 6
rect 550 -97 1198 -93
rect 1201 -2 1230 2
rect 1201 -102 1205 -2
rect 541 -106 1205 -102
rect 1208 -10 1229 -6
rect 1208 -111 1212 -10
rect 532 -115 1212 -111
rect 1215 -18 1231 -14
rect 1215 -120 1219 -18
rect 523 -124 1219 -120
<< m2contact >>
rect 505 177 510 182
rect 917 54 922 59
rect 544 31 549 36
rect 1225 54 1230 59
rect 535 23 540 28
rect 526 15 531 20
rect 517 7 522 12
rect 504 -49 509 -44
rect 545 -97 550 -92
rect 536 -106 541 -101
rect 527 -115 532 -110
rect 518 -124 523 -119
<< metal2 >>
rect 505 -44 509 177
rect 922 54 1225 58
rect 518 -119 522 7
rect 527 -110 531 15
rect 536 -101 540 23
rect 545 -92 549 31
use PG  PG_0
timestamp 1638826306
transform 1 0 39 0 1 82
box -39 -152 461 111
use CLA  CLA_0
timestamp 1638826311
transform 1 0 613 0 1 58
box -41 -147 565 328
use SUM  SUM_0
timestamp 1638824961
transform 1 0 1254 0 1 54
box -28 -72 485 109
<< end >>
