* SPICE3 file created from and3.ext - technology: scmos

.option scale=0.09u

M1000 out nandout vdd w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=152 ps=86
M1001 nandout C a_24_n25# Gnd nfet w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1002 vdd B nandout w_0_0# pfet w=8 l=2
+  ad=0 pd=0 as=112 ps=60
M1003 a_24_n25# B a_14_n25# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1004 a_14_n25# A gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=44 ps=38
M1005 nandout A vdd w_0_0# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 nandout C vdd w_0_0# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 out nandout gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
