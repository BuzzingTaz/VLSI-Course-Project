* SPICE3 file created from SUM.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY=1.8
.option scale=0.09u
.global vdd gnd

Vdd vdd gnd SUPPLY
vA0 P0 gnd pulse 0 1.8 0us 100ps 100ps 9.9us 20us
vA1 P1 gnd pulse 0 1.8 0us 100ps 100ps 9.9us 20us
vA2 P2 gnd pulse 0 1.8 0us 100ps 100ps 9.9us 20us
vA3 P3 gnd pulse 0 1.8 0us 100ps 100ps 9.9us 20us
vB0 C4 gnd pulse 0 1.8 0us 100ps 100ps 19.8us 40us
vB1 C1 gnd pulse 0 1.8 0us 100ps 100ps 19.8us 40us
vB2 C2 gnd pulse 0 1.8 0us 100ps 100ps 19.8us 40us
vB3 C3 gnd pulse 0 1.8 0us 100ps 100ps 19.8us 40us
vC0 C0 gnd pulse 0 1.8 0us 100ps 100ps 19.6us 40us

M1000 xor_0/Bbar C0 vdd xor_0/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=640 ps=352
M1001 xor_0/Bbar C0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=384 ps=320
M1002 S0 C0 xor_0/a_15_n48# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1003 vdd P0 xor_0/a_7_6# xor_0/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=160 ps=88
M1004 xor_0/a_15_n48# P0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 xor_0/Abar P0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1006 xor_0/a_7_6# xor_0/Bbar S0 xor_0/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1007 S0 xor_0/Abar xor_0/a_7_6# xor_0/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 xor_0/Abar P0 vdd xor_0/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1009 gnd xor_0/Bbar xor_0/a_35_n48# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1010 xor_0/a_7_6# C0 vdd xor_0/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 xor_0/a_35_n48# xor_0/Abar S0 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 xor_1/Bbar C1 vdd xor_1/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1013 xor_1/Bbar C1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1014 S1 C1 xor_1/a_15_n48# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1015 vdd P1 xor_1/a_7_6# xor_1/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=160 ps=88
M1016 xor_1/a_15_n48# P1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 xor_1/Abar P1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1018 xor_1/a_7_6# xor_1/Bbar S1 xor_1/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1019 S1 xor_1/Abar xor_1/a_7_6# xor_1/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 xor_1/Abar P1 vdd xor_1/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1021 gnd xor_1/Bbar xor_1/a_35_n48# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1022 xor_1/a_7_6# C1 vdd xor_1/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 xor_1/a_35_n48# xor_1/Abar S1 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 xor_2/Bbar C2 vdd xor_2/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1025 xor_2/Bbar C2 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1026 S2 C2 xor_2/a_15_n48# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1027 vdd P2 xor_2/a_7_6# xor_2/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=160 ps=88
M1028 xor_2/a_15_n48# P2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 xor_2/Abar P2 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1030 xor_2/a_7_6# xor_2/Bbar S2 xor_2/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1031 S2 xor_2/Abar xor_2/a_7_6# xor_2/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 xor_2/Abar P2 vdd xor_2/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1033 gnd xor_2/Bbar xor_2/a_35_n48# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1034 xor_2/a_7_6# C2 vdd xor_2/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 xor_2/a_35_n48# xor_2/Abar S2 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 xor_3/Bbar C3 vdd xor_3/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1037 xor_3/Bbar C3 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1038 S3 C3 xor_3/a_15_n48# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1039 vdd P3 xor_3/a_7_6# xor_3/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=160 ps=88
M1040 xor_3/a_15_n48# P3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 xor_3/Abar P3 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1042 xor_3/a_7_6# xor_3/Bbar S3 xor_3/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1043 S3 xor_3/Abar xor_3/a_7_6# xor_3/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 xor_3/Abar P3 vdd xor_3/w_n35_0# CMOSP w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1045 gnd xor_3/Bbar xor_3/a_35_n48# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1046 xor_3/a_7_6# C3 vdd xor_3/w_n35_0# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 xor_3/a_35_n48# xor_3/Abar S3 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 P3 P2 2.68fF
C1 C3 C2 2.77fF
C2 gnd Gnd 2.79fF
C3 vdd Gnd 2.73fF
C4 P3 Gnd 2.93fF
C5 C3 Gnd 3.22fF
C6 P2 Gnd 2.46fF
C7 C2 Gnd 2.71fF
C8 C1 Gnd 2.19fF


.tran 10n 80us

.control
run

plot v(P0)

plot v(P1)

plot v(P2)
plot  v(P3)

plot v(S0)
plot v(S1)
plot v(S2)
plot v(S3)

.endc
.end