magic
tech scmos
timestamp 1638771050
<< nwell >>
rect 0 3 61 23
<< ntransistor >>
rect 11 -22 13 -18
rect 21 -22 23 -18
rect 31 -22 33 -18
rect 48 -22 50 -18
<< ptransistor >>
rect 11 9 13 17
rect 21 9 23 17
rect 31 9 33 17
rect 48 9 50 17
<< ndiffusion >>
rect 10 -22 11 -18
rect 13 -22 15 -18
rect 19 -22 21 -18
rect 23 -22 25 -18
rect 29 -22 31 -18
rect 33 -22 35 -18
rect 47 -22 48 -18
rect 50 -22 51 -18
<< pdiffusion >>
rect 10 9 11 17
rect 13 9 21 17
rect 23 9 31 17
rect 33 9 35 17
rect 47 9 48 17
rect 50 9 51 17
<< ndcontact >>
rect 6 -22 10 -18
rect 15 -22 19 -18
rect 25 -22 29 -18
rect 35 -22 39 -18
rect 43 -22 47 -18
rect 51 -22 55 -18
<< pdcontact >>
rect 6 9 10 17
rect 35 9 39 17
rect 43 9 47 17
rect 51 9 55 17
<< polysilicon >>
rect 11 17 13 20
rect 21 17 23 20
rect 31 17 33 20
rect 48 17 50 20
rect 11 -18 13 9
rect 21 -18 23 9
rect 31 -18 33 9
rect 48 -18 50 9
rect 11 -25 13 -22
rect 21 -25 23 -22
rect 31 -25 33 -22
rect 48 -25 50 -22
<< polycontact >>
rect 7 -15 11 -11
rect 17 -8 21 -4
rect 27 -1 31 3
rect 44 -15 48 -11
<< metal1 >>
rect 0 23 61 27
rect 6 17 10 23
rect 43 17 47 23
rect 0 -1 27 3
rect 0 -8 17 -4
rect 35 -11 39 9
rect 51 -7 55 9
rect 51 -11 61 -7
rect 0 -15 7 -11
rect 15 -15 44 -11
rect 15 -18 19 -15
rect 35 -18 39 -15
rect 51 -18 55 -11
rect 6 -26 10 -22
rect 25 -26 29 -22
rect 43 -26 47 -22
rect 0 -30 61 -26
<< labels >>
rlabel metal1 1 25 1 25 4 vdd
rlabel metal1 29 25 29 25 4 vdd
rlabel metal1 1 -28 1 -28 2 gnd
rlabel metal1 57 -9 57 -9 7 orout
rlabel metal1 2 1 2 1 3 C
rlabel metal1 2 -6 2 -6 3 B
rlabel metal1 2 -13 2 -13 3 A
<< end >>
