magic
tech scmos
timestamp 1638782314
<< nwell >>
rect 0 3 71 23
<< ntransistor >>
rect 11 -29 13 -25
rect 21 -29 23 -25
rect 31 -29 33 -25
rect 41 -29 43 -25
rect 58 -29 60 -25
<< ptransistor >>
rect 11 9 13 17
rect 21 9 23 17
rect 31 9 33 17
rect 41 9 43 17
rect 58 9 60 17
<< ndiffusion >>
rect 10 -29 11 -25
rect 13 -29 15 -25
rect 19 -29 21 -25
rect 23 -29 25 -25
rect 29 -29 31 -25
rect 33 -29 41 -25
rect 43 -29 45 -25
rect 57 -29 58 -25
rect 60 -29 61 -25
<< pdiffusion >>
rect 10 9 11 17
rect 13 9 21 17
rect 23 9 31 17
rect 33 9 41 17
rect 43 9 45 17
rect 57 9 58 17
rect 60 9 61 17
<< ndcontact >>
rect 6 -29 10 -25
rect 15 -29 19 -25
rect 25 -29 29 -25
rect 45 -29 49 -25
rect 53 -29 57 -25
rect 61 -29 65 -25
<< pdcontact >>
rect 6 9 10 17
rect 45 9 49 17
rect 53 9 57 17
rect 61 9 65 17
<< polysilicon >>
rect 11 17 13 20
rect 21 17 23 20
rect 31 17 33 20
rect 41 17 43 20
rect 58 17 60 20
rect 11 -25 13 9
rect 21 -25 23 9
rect 31 -25 33 9
rect 41 -25 43 9
rect 58 -25 60 9
rect 11 -32 13 -29
rect 21 -32 23 -29
rect 31 -32 33 -29
rect 41 -32 43 -29
rect 58 -32 60 -29
<< polycontact >>
rect 7 -22 11 -18
rect 17 -15 21 -11
rect 27 -8 31 -4
rect 37 -1 41 3
rect 54 -22 58 -18
<< metal1 >>
rect 0 23 71 27
rect 6 17 10 23
rect 53 17 57 23
rect 0 -1 37 3
rect 0 -8 27 -4
rect 0 -15 17 -11
rect 45 -18 49 9
rect 61 3 65 9
rect 61 -1 71 3
rect 0 -22 7 -18
rect 15 -22 54 -18
rect 15 -25 19 -22
rect 35 -29 39 -22
rect 61 -25 65 -1
rect 6 -33 10 -29
rect 25 -33 29 -29
rect 45 -33 49 -29
rect 53 -33 57 -29
rect 0 -37 71 -33
<< labels >>
rlabel metal1 1 25 1 25 4 vdd
rlabel metal1 29 25 29 25 4 vdd
rlabel metal1 1 1 1 1 3 D
rlabel metal1 1 -35 1 -35 2 gnd
rlabel metal1 2 -6 2 -6 3 C
rlabel metal1 2 -13 2 -13 3 B
rlabel metal1 2 -20 2 -20 3 A
rlabel metal1 67 1 67 1 7 orout
<< end >>
