magic
tech scmos
timestamp 1638829229
<< metal1 >>
rect 1172 382 1230 386
rect 1177 351 1212 355
rect 495 238 583 242
rect 495 169 499 238
rect 1037 214 1213 218
rect 510 178 586 182
rect -4 165 0 169
rect 485 165 499 169
rect -4 82 0 86
rect 924 82 1206 83
rect 921 79 1206 82
rect -4 74 0 78
rect -4 67 0 71
rect -4 60 0 64
rect 917 59 921 64
rect -4 53 0 57
rect -4 45 0 49
rect 498 45 576 49
rect -4 37 0 41
rect 1202 39 1206 79
rect 1209 47 1213 214
rect 1226 137 1230 382
rect 1244 351 1740 355
rect 1736 135 1740 351
rect 1736 131 1743 135
rect 1739 119 1743 123
rect 1739 111 1743 115
rect 1739 103 1743 107
rect 1739 91 1743 95
rect 1209 43 1230 47
rect -4 30 0 34
rect 498 31 517 35
rect 1202 35 1227 39
rect 1229 35 1232 39
rect 522 31 576 35
rect -4 23 0 27
rect 497 23 526 27
rect 1187 27 1230 31
rect 531 23 575 27
rect -4 16 0 20
rect 499 15 535 19
rect 540 15 577 19
rect 499 7 544 11
rect 549 7 577 11
rect 486 -2 576 2
rect 483 -11 576 -7
rect 484 -20 577 -16
rect 485 -27 578 -23
rect 496 -49 504 -45
rect 1187 -63 1191 27
rect 828 -66 1191 -63
rect 831 -67 1191 -66
rect 1194 6 1234 10
rect 1194 -93 1198 6
rect 550 -97 1198 -93
rect 1201 -2 1230 2
rect 1201 -102 1205 -2
rect 541 -106 1205 -102
rect 1208 -10 1229 -6
rect 1208 -111 1212 -10
rect 532 -115 1212 -111
rect 1215 -18 1231 -14
rect 1215 -120 1219 -18
rect 523 -124 1219 -120
<< m2contact >>
rect 1212 351 1217 356
rect 505 177 510 182
rect 917 54 922 59
rect 937 44 942 49
rect 1239 351 1244 356
rect 1225 54 1230 59
rect 517 31 522 36
rect 526 23 531 28
rect 535 15 540 20
rect 544 6 549 11
rect 504 -49 509 -44
rect 1226 18 1231 23
rect 545 -97 550 -92
rect 536 -106 541 -101
rect 527 -115 532 -110
rect 518 -124 523 -119
<< metal2 >>
rect 1217 351 1239 355
rect 505 -44 509 177
rect 922 54 1225 58
rect 518 -119 522 31
rect 527 -110 531 23
rect 938 23 942 44
rect 938 19 1226 23
rect 536 -101 540 15
rect 545 -92 549 6
use PG  PG_0
timestamp 1638826306
transform 1 0 39 0 1 82
box -39 -152 461 111
use CLA  CLA_0
timestamp 1638828401
transform 1 0 613 0 1 58
box -41 -147 565 328
use SUM  SUM_0
timestamp 1638824961
transform 1 0 1254 0 1 54
box -28 -72 485 109
<< labels >>
rlabel metal1 1741 93 1741 93 7 S0
rlabel metal1 1741 105 1741 105 7 S1
rlabel metal1 1741 113 1741 113 7 S2
rlabel metal1 1741 121 1741 121 7 S3
rlabel metal1 1741 133 1741 133 7 Cout
rlabel metal1 -2 84 -2 84 3 gnd
rlabel metal1 -2 76 -2 76 3 A0
rlabel metal1 -2 69 -2 69 3 A1
rlabel metal1 -2 62 -2 62 3 A2
rlabel metal1 -2 55 -2 55 3 A3
rlabel metal1 -2 47 -2 47 3 C0
rlabel metal1 -2 39 -2 39 3 B0
rlabel metal1 -2 32 -2 32 3 B1
rlabel metal1 -2 25 -2 25 3 B2
rlabel metal1 -2 18 -2 18 3 B3
<< end >>
