magic
tech scmos
timestamp 1638780161
<< nwell >>
rect 0 3 50 23
<< ntransistor >>
rect 11 -15 13 -11
rect 21 -15 23 -11
rect 37 -15 39 -11
<< ptransistor >>
rect 11 9 13 17
rect 21 9 23 17
rect 37 9 39 17
<< ndiffusion >>
rect 10 -15 11 -11
rect 13 -15 21 -11
rect 23 -15 24 -11
rect 36 -15 37 -11
rect 39 -15 40 -11
<< pdiffusion >>
rect 10 9 11 17
rect 13 9 15 17
rect 19 9 21 17
rect 23 9 24 17
rect 36 9 37 17
rect 39 9 40 17
<< ndcontact >>
rect 6 -15 10 -11
rect 24 -15 28 -11
rect 32 -15 36 -11
rect 40 -15 44 -11
<< pdcontact >>
rect 6 9 10 17
rect 15 9 19 17
rect 24 9 28 17
rect 32 9 36 17
rect 40 9 44 17
<< polysilicon >>
rect 11 17 13 20
rect 21 17 23 20
rect 37 17 39 20
rect 11 -11 13 9
rect 21 -11 23 9
rect 37 -11 39 9
rect 11 -18 13 -15
rect 21 -18 23 -15
rect 37 -18 39 -15
<< polycontact >>
rect 7 -1 11 3
rect 17 -8 21 -4
rect 33 -1 37 3
<< metal1 >>
rect 0 23 50 27
rect 6 17 10 23
rect 24 17 28 23
rect 32 17 36 23
rect 15 3 19 9
rect 40 3 44 9
rect 0 -1 7 3
rect 15 -1 33 3
rect 40 -1 50 3
rect 0 -8 17 -4
rect 24 -11 28 -1
rect 40 -11 44 -1
rect 6 -19 10 -15
rect 32 -19 36 -15
rect 0 -23 50 -19
<< labels >>
rlabel metal1 1 25 1 25 4 vdd
rlabel metal1 16 -6 16 -6 1 B
rlabel metal1 6 1 6 1 1 A
rlabel metal1 1 -21 1 -21 2 gnd
rlabel metal1 46 0 46 0 7 andout
<< end >>
