magic
tech scmos
timestamp 1638800402
<< nwell >>
rect 0 3 81 23
<< ntransistor >>
rect 11 -36 13 -32
rect 21 -36 23 -32
rect 31 -36 33 -32
rect 41 -36 43 -32
rect 51 -36 53 -32
rect 68 -36 70 -32
<< ptransistor >>
rect 11 9 13 17
rect 21 9 23 17
rect 31 9 33 17
rect 41 9 43 17
rect 51 9 53 17
rect 68 9 70 17
<< ndiffusion >>
rect 10 -36 11 -32
rect 13 -36 15 -32
rect 19 -36 21 -32
rect 23 -36 25 -32
rect 29 -36 31 -32
rect 33 -36 41 -32
rect 43 -36 45 -32
rect 49 -36 51 -32
rect 53 -36 55 -32
rect 67 -36 68 -32
rect 70 -36 71 -32
<< pdiffusion >>
rect 10 9 11 17
rect 13 9 21 17
rect 23 9 31 17
rect 33 9 41 17
rect 43 9 51 17
rect 53 9 55 17
rect 67 9 68 17
rect 70 9 71 17
<< ndcontact >>
rect 6 -36 10 -32
rect 15 -36 19 -32
rect 25 -36 29 -32
rect 45 -36 49 -32
rect 55 -36 59 -32
rect 63 -36 67 -32
rect 71 -36 75 -32
<< pdcontact >>
rect 6 9 10 17
rect 55 9 59 17
rect 63 9 67 17
rect 71 9 75 17
<< polysilicon >>
rect 11 17 13 20
rect 21 17 23 20
rect 31 17 33 20
rect 41 17 43 20
rect 51 17 53 20
rect 68 17 70 20
rect 11 -32 13 9
rect 21 -32 23 9
rect 31 -32 33 9
rect 41 -32 43 9
rect 51 -32 53 9
rect 68 -32 70 9
rect 11 -39 13 -36
rect 21 -39 23 -36
rect 31 -39 33 -36
rect 41 -39 43 -36
rect 51 -39 53 -36
rect 68 -39 70 -36
<< polycontact >>
rect 7 -29 11 -25
rect 17 -22 21 -18
rect 27 -15 31 -11
rect 37 -8 41 -4
rect 47 -1 51 3
rect 64 -29 68 -25
<< metal1 >>
rect 0 23 81 27
rect 6 17 10 23
rect 63 17 67 23
rect 0 -1 47 3
rect 0 -8 37 -4
rect 0 -15 27 -11
rect 0 -22 17 -18
rect 55 -25 59 9
rect 71 -4 75 9
rect 71 -8 81 -4
rect 0 -29 7 -25
rect 15 -29 64 -25
rect 15 -32 19 -29
rect 35 -36 39 -29
rect 55 -32 59 -29
rect 71 -32 75 -8
rect 6 -40 10 -36
rect 25 -40 29 -36
rect 45 -40 49 -36
rect 63 -40 67 -36
rect 0 -44 81 -40
<< labels >>
rlabel metal1 1 25 1 25 4 vdd
rlabel metal1 29 25 29 25 4 vdd
rlabel metal1 1 -6 1 -6 3 D
rlabel metal1 1 -42 1 -42 2 gnd
rlabel metal1 2 -13 2 -13 3 C
rlabel metal1 2 -20 2 -20 3 B
rlabel metal1 2 -27 2 -27 3 A
rlabel metal1 77 -6 77 -6 7 orout
rlabel metal1 1 1 1 1 3 E
<< end >>
