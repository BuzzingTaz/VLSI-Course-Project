magic
tech scmos
timestamp 1638797340
<< nwell >>
rect 0 0 82 20
<< ntransistor >>
rect 12 -39 14 -35
rect 22 -39 24 -35
rect 32 -39 34 -35
rect 42 -39 44 -35
rect 52 -39 54 -35
rect 69 -39 71 -35
<< ptransistor >>
rect 12 6 14 14
rect 22 6 24 14
rect 32 6 34 14
rect 42 6 44 14
rect 52 6 54 14
rect 69 6 71 14
<< ndiffusion >>
rect 10 -39 12 -35
rect 14 -39 22 -35
rect 24 -39 32 -35
rect 34 -39 42 -35
rect 44 -39 52 -35
rect 54 -39 56 -35
rect 68 -39 69 -35
rect 71 -39 72 -35
<< pdiffusion >>
rect 10 6 12 14
rect 14 6 16 14
rect 20 6 22 14
rect 24 6 26 14
rect 30 6 32 14
rect 34 6 36 14
rect 40 6 42 14
rect 44 6 46 14
rect 50 6 52 14
rect 54 6 56 14
rect 68 6 69 14
rect 71 6 72 14
<< ndcontact >>
rect 6 -39 10 -35
rect 56 -39 60 -35
rect 64 -39 68 -35
rect 72 -39 76 -35
<< pdcontact >>
rect 6 6 10 14
rect 16 6 20 14
rect 26 6 30 14
rect 36 6 40 14
rect 46 6 50 14
rect 56 6 60 14
rect 64 6 68 14
rect 72 6 76 14
<< polysilicon >>
rect 12 14 14 17
rect 22 14 24 17
rect 32 14 34 17
rect 42 14 44 17
rect 52 14 54 17
rect 69 14 71 17
rect 12 -35 14 6
rect 22 -35 24 6
rect 32 -35 34 6
rect 42 -35 44 6
rect 52 -35 54 6
rect 69 -35 71 6
rect 12 -42 14 -39
rect 22 -42 24 -39
rect 32 -42 34 -39
rect 42 -42 44 -39
rect 52 -42 54 -39
rect 69 -42 71 -39
<< polycontact >>
rect 8 -4 12 0
rect 18 -11 22 -7
rect 28 -18 32 -14
rect 38 -25 42 -21
rect 48 -32 52 -28
rect 65 -4 69 0
<< metal1 >>
rect 0 20 82 24
rect 6 14 10 20
rect 26 14 30 20
rect 46 14 50 20
rect 64 14 68 20
rect 16 0 20 6
rect 36 0 40 6
rect 56 0 60 6
rect 72 0 76 6
rect 0 -4 8 0
rect 16 -4 65 0
rect 72 -4 82 0
rect 0 -11 18 -7
rect 0 -18 28 -14
rect 0 -25 38 -21
rect 0 -32 48 -28
rect 56 -35 60 -4
rect 72 -35 76 -4
rect 6 -43 10 -39
rect 64 -43 68 -39
rect 0 -47 82 -43
<< labels >>
rlabel metal1 1 -9 1 -9 3 B
rlabel metal1 2 22 2 22 4 vdd
rlabel metal1 1 -23 1 -23 3 D
rlabel metal1 1 -16 1 -16 3 C
rlabel metal1 1 -2 1 -2 3 A
rlabel metal1 80 -2 80 -2 7 out
rlabel metal1 2 -45 2 -45 2 gnd
rlabel metal1 1 -30 1 -30 3 E
<< end >>
